// TIMESTAMP.vh
// Sun Sep 25 12:06:52 JST 2022
// 632FC5CC
parameter [31:0] C_TIMESTAMP = 32'h632FC5CC ;
