`include "./TIMESTAMP.vh"
// {C_USEs[7:0],C_DEFAULTs[7:0]} //1address
parameter C_INITss = {
    {256{8'b0000_0000,8'b0000_0000}}
    ,{8'b0000_0000,8'b0000_0000}    //0F
    ,{8'b0000_0000,8'b0000_0000}    //0E
    ,{8'b0000_0000,8'b0000_0000}    //0D
    ,{8'b0000_0000,8'b0000_0000}    //0C
    ,{8'b0000_0000,8'b0000_0000}    //0B
    ,{8'b0000_0000,8'b0000_0000}    //0A
    ,{8'b1111_1111,8'b1111_0000}    //09
    ,{8'b1111_1111,8'b1010_0101}    //08    //                              
    ,{8'b0000_0000,C_TIMESTAMP[3*8+:8]} //07 version
    ,{8'b0000_0000,C_TIMESTAMP[2*8+:8]} //06
    ,{8'b0000_0000,C_TIMESTAMP[1*8+:8]} //05
    ,{8'b0000_0000,C_TIMESTAMP[0*8+:8]} //04
    ,{8'b0000_0000,8'h76}               //03 time_stamp
    ,{8'b0000_0000,8'h54}               //02
    ,{8'b0000_0000,8'h32}               //01
    ,{8'b0000_0000,8'h10}               //00
};
