// TIMESTAMP.vh
// Sun Sep 25 18:38:18 JST 2022
// 6330218A
parameter [31:0] C_TIMESTAMP = 32'h6330218A ;
