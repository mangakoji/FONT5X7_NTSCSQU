// TIMESTAMP.vh
// Sun Sep 25 21:29:56 JST 2022
// 633049C4
parameter [31:0] C_TIMESTAMP = 32'h633049C4 ;
